module Top
(
);

endmodule