module ADC_Interface
(
    output CLKOUT,
    input MISO[11:0]
);

endmodule